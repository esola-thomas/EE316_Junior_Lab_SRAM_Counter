ROM_inst : ROM PORT MAP (
		address	 => address_sig,
		clken	 => clken_sig,
		clock	 => clock_sig,
		q	 => q_sig
	);
